class abc;
  rand int a[];
  
  constraint c1{a.size==100;}
  
  constraint c3{foreach(a[i]) if(i<4) a[i]==i+1;
                else if(i>=4) 
  						{
                  if(i%4==0) a[i] == a[i-4]+1;
                  else if(i%4==1) a[i] == a[i-4]+1;
                  else if(i%4==2) a[i] == a[i-4]+1;
                  else if(i%4==3) a[i] == a[i-4]+1;
                }
               }

endclass

module m1;
  
  abc p;
  
  initial begin
    p = new();
    
    p.randomize();
    $display("a[]=%p",p.a);
  end
endmodule


------------------------------------------------------------------------------------------------------------------------------------
                              V C S   S i m u l a t i o n   R e p o r t
------------------------------------------------------------------------------------------------------------------------------------
a[]='{1, 2, 3, 4, 2, 3, 4, 5, 3, 4, 5, 6, 4, 5, 6, 7, 5, 6, 7, 8, 6, 7, 8, 9, 7, 8, 9, 10, 8, 9, 10, 11, 9, 10, 11, 12, 10, 11, 12, 
      13, 11, 12, 13, 14, 12, 13, 14, 15, 13, 14, 15, 16, 14, 15, 16, 17, 15, 16, 17, 18, 16, 17, 18, 19, 17, 18, 19, 20, 18, 19, 20, 
      21, 19, 20, 21, 22, 20, 21, 22, 23, 21, 22, 23, 24, 22, 23, 24, 25, 23, 24, 25, 26, 24, 25, 26, 27, 25, 26, 27, 28} 
------------------------------------------------------------------------------------------------------------------------------------
