class A;
  rand logic [31:0] a;
  int i;
  constraint C1 { foreach(a[i]) 
                    if(i%2 ==0) 
                      a[i] == 0;
                 	  else 
                   	  a[i] == 1;
                }
endclass
  
module test;        
  A a1;
    
  initial begin 
     a1 = new();
     repeat(10)
      begin
        a1.randomize();
        $display(" a = %0b",a1.a);
      end 
  end 
endmodule

-------------------------------------------------------------------------------------
                 V C S   S i m u l a t i o n   R e p o r t
-------------------------------------------------------------------------------------

 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
 a = 10101010101010101010101010101010
-------------------------------------------------------------------------------------
