class prime;
  rand int q[$];
  constraint c1{ q.size inside {[30:100]};
                    foreach(q[i])
                      if(((i%2==0 && i!=2) || (i%3==0 && i!=3)  || (i%4==0 && i!=4) || (i%5==0 && i!=5) || (i%6==0 && i!=6) || (i%7==0 && i!=7) || (i%8==0 && i!=8) || (i%9==0 && i!=9)))

                         q[i]==1;
                      else
                        q[i]==i; }

  function void disp();
    $display("q: %p",q);
  endfunction
endclass

module m1;
  prime a1;
  initial begin
    a1=new();
    a1.randomize();
    a1.disp();
  end
endmodule


---------------------------------------------------------------------------------------------------------------------------------------------------
                                           V C S   S i m u l a t i o n   R e p o r t 
---------------------------------------------------------------------------------------------------------------------------------------------------
q: '{1, 1, 2, 3, 1, 5, 1, 7, 1, 1, 1, 11, 1, 13, 1, 1, 1, 17, 1, 19, 1, 1, 1, 23, 1, 1, 1, 1, 1, 29, 1, 31, 1, 1, 1, 1, 1, 37, 1, 1, 1, 41, 1, 43}
---------------------------------------------------------------------------------------------------------------------------------------------------
